LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use work.mypack.all;

ENTITY tb_MulUnit IS
END tb_MulUnit;
 
ARCHITECTURE behavior OF tb_MulUnit IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT MultiplierUnit_7x7_to_49
    PORT(
         image : IN  matrix;
         coefficient : IN  matrix;
         result : OUT  line
        );
    END COMPONENT;
    

   --Inputs
   signal image : matrix;
   signal coefficient : matrix;

 	--Outputs
   signal result : line;

  
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: MultiplierUnit_7x7_to_49 PORT MAP (
          image => image,
          coefficient => coefficient,
          result => result
        );


   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		image <= ((("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")));
		
		coefficient <= ((("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")),
		(("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010"),("00000010")));
      -- insert stimulus here 

      wait;
   end process;

END;
